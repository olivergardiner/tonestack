Tube Driver circuit for tonestack

* Insert you circuit in the area marked below - do not change anything else.
* The input to your circuit is node 2 relative to node 0 which is ground
* The output of your circuit must be node 3

* Four potentiometers are nominally available for you to use in your circuit:
* Pot 1 must consist of RP1LO and RP1HI
* Pot 2 must consist of RP2LO and RP2HI
* Pot 3 must consist of RP3LO and RP3HI
* Pot 4 must consist of RP4LO and RP4HI - this is currently inactive

* Nodes 0 to 9 are reserved

VIN 0 1 DC 0 AC 1
R98 1 2 38K

******* PLACE YOUR CIRCUIT HERE *******

R1 2 10 22K
C1 2 11 330P
C2 10 12 100N
C3 10 13 47N
R2 13 0 22K
C4 13 0 47N
R3 3 12 220K

RP1LO 13 12 10K
RP1HI 12 12 90K

RP3LO 12 3 50K
RP3HI 3 11 450K

******* PLACE YOUR CIRCUIT HERE *******

R99 3 0 100K

.OPTIONS NOACCT
.AC DEC 40 10 100K

.END