Vortex Drive filter circuit for tonestack

* Insert you circuit in the area marked below - do not change anything else.
* The input to your circuit is node 2 relative to node 0 which is ground
* The output of your circuit must be node 3

* Four potentiometers are nominally available for you to use in your circuit:
* Pot 1 must consist of RP1LO and RP1HI
* Pot 2 must consist of RP2LO and RP2HI
* Pot 3 must consist of RP3LO and RP3HI
* Pot 4 must consist of RP4LO and RP4HI - this is cuurently inactive

* Nodes 0 to 9 are reserved

VIN 0 1 DC 0 AC 1
R98 1 2 47

******* PLACE YOUR CIRCUIT HERE *******
.INCLUDE OPAMP1.cir

R1 13 15 200K
R2 16 0  8.2K
R3 12 18 470K
C1 12 14 4.7N
C2 13 14 4.7N
C3 18 13 4.7N

RP1LO 3 10 8K
RP1HI 10 2 2K

RP3LO 15 16 70K
RP3HI 16 14 30K

XOPAMP1 10 12 18 OPAMP1

RD1 18 21 22K
RD2 10 20 22K
RD3 21 0 22K
RD4 20 22 22K
XOPAMP2 21 20 22 OPAMP1

RS1 2 30 10K
RS2 22 30 10K
RS3 30 3 10K
XOPAMP3 0 30 3 OPAMP1

******* PLACE YOUR CIRCUIT HERE *******

R99 3 0 10K

.OPTIONS NOACCT
.AC DEC 40 10 100K

.END