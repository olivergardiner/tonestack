Vox circuit for tonestack

* Insert you circuit in the area marked below - do not change anything else.
* The input to your circuit is node 2 relative to node 0 which is ground
* The output of your circuit must be node 3

* Four potentiometers are nominally available for you to use in your circuit:
* Pot 1 must consist of RP1LO and RP1HI
* Pot 2 must consist of RP2LO and RP2HI
* Pot 3 must consist of RP3LO and RP3HI
* Pot 4 must consist of RP4LO and RP4HI - this is currently inactive

* Nodes 0 to 9 are reserved

VIN 0 1 DC 0 AC 1
R98 1 2 56K

******* PLACE YOUR CIRCUIT HERE *******

R1 2 10 100K
C1 10 12 22N
C2 10 13 22N
C3 2 11 47P
R2 12 0 10K

* Bass 1M LogA
RP1LO 12 13 500K
RP1HI 0 12 500K

* Treble 1M Log A
RP3LO 13 3 500K
RP3HI 3 11 500K

******* PLACE YOUR CIRCUIT HERE *******

R99 3 0 1MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END