* OPAMP2.CIR - OPAMP MODEL (LEVEL 2)
* OPAMP MACRO MODEL (INTERMEDIATE LEVEL)
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | |   NEGATIVE POWER SUPPLY
*                | | |   |   OUTPUT
*                | | |   |   |
.SUBCKT OPAMP2   1 2 101 102 81  
Q1	5 1	7	NPN
Q2	6 2	8	NPN
RC1	101	5	95.49
RC2	101	6	95.49
RE1	7	4	43.79
RE2	8	4	43.79
I1	4	102	0.001
*
* OPEN-LOOP GAIN, FIRST POLE AND SLEW RATE
G1	100 10	6 5 0.0104719
RP1	10	100	9.549MEG
CP1	10	100	0.0016667UF
*
*OUTPUT STAGE
EOUT	80 100	10 100	1
RO	80	81	100
*
* INTERNAL REFERENCE
RREF1	101	103	100K
RREF2	103	102	100K
EREF	100 0	103 0 1
R100	100	0	1MEG
*
.model NPN  NPN(BF=50000)
*
.ENDS