Single control tone circuit #1

VIN 0 1 DC 0 AC 1
RS 1 2 47K

R1 2 4 220K

RTONEHI 4 5 250K
RTONELO 5 0 250K

R2 2 6 470K
C1 5 6 560p
R3 6 0 270K

RVOLHI 6 3 1
RVOLLO 3 0 1MEG

RL 3 0 10MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END