Vortex Drive filter circuit for tonestack

* Insert you circuit in the area marked below - do not change anything else.
* The input to your circuit is node 2 relative to node 0 which is ground
* The output of your circuit must be node 3

* Four potentiometers are nominally available for you to use in your circuit:
* Pot 1 must consist of RP1LO and RP1HI
* Pot 2 must consist of RP2LO and RP2HI
* Pot 3 must consist of RP3LO and RP3HI
* Pot 4 must consist of RP4LO and RP4HI - this is currently inactive

* Nodes 0 to 9 are reserved

VIN 0 1 DC 0 AC 1
R98 1 2 820

******* PLACE YOUR CIRCUIT HERE *******
.INCLUDE OPAMP1.cir

.MODEL 2SC1815 NPN (IS=9.99315F BF=192.019 NF=1.01109 VAF=311.281 IKF=214.789M
+ ISE=124.464F NE=1.51791 BR=4.99998 IKR=980.183 ISC=33.4247F RE=2.96389 CJE=2P
+ MJE=500M CJC=7.82341P VJC=700M MJC=500.188M TF=512.206P XTF=183.171M
+ VTF=9.97698 ITF=9.76409M TR=10N )

.MODEL NPN NPN

VCC 0 40 DC 9
VB  0 41 DC 4.5

R1 2  10 9.1K
R2 10 11 10K
R3 12 13 39K
R4 12 3  82K
R5 16 19 1K

C1 2  0  100N
C2 11 0  10N
C3 13 0  100N
C4 15 16 33N
C5 16 17 10N

RLIM  12 18 100R
RP2HI 18 15 50K
RP2LO 15 14 50K

XOPAMP1 11 12 3  OPAMP1
* CX 12 3  47P

Q1 40 17 19 2SC1815
RE 19 0  10K
RB 17 41 100K

* XOPAMP2 17 19 19 OPAMP1

******* PLACE YOUR CIRCUIT HERE *******

R99 3 0 10K

.OPTIONS NOACCT
.AC DEC 40 10 100K

.END