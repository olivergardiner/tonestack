Fender classic three knob control

VIN 0 1 DC 0 AC 1
RS 1 2 56K

C1 2 4 47P
R1 2 5 100K

RTREBLEHI 4 7 500K
RTREBLELO 7 6 500K

C2 5 6 22N
C3 5 9 22N
R2 9 0 10K

RBASSHI 6 9 500K
RBASSLO 0 9 500K

RVOLHI 7 3 1
RVOLLO 3 0 600K

RL 3 0 10MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END