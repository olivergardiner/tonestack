* OPMODEL1.CIR - OPAMP MODEL SINGLE-POLE
* OPAMP MACRO MODEL (BASIC LEVEL)
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | OUTPUT
*                | | |
.SUBCKT OPAMP1	 1 2 6
* INPUT IMPEDANCE
RIN	1	2	10MEG
* DC GAIN=100K AND POLE1=100HZ
* UNITY GAIN = DCGAIN X POLE1 = 10MHZ
EGAIN	3 0	1 2	100K
RP1	3	4	1K
CP1	4	0	1.5915UF
* OUTPUT BUFFER AND RESISTANCE
EBUFFER	5 0	4 0	1
ROUT	5	6	10
.ENDS