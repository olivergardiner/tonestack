Marshall classic three knob control

VIN 0 1 DC 0 AC 1
RS 1 2 1

C1 2 4 470P
R1 2 5 33K

RTREBLEHI 4 7 110K
RTREBLELO 7 6 110K

C2 5 6 22N
C3 5 8 22N

RMIDHI 9 8 12.5K
RMIDLO 8 0 12.5K

RBASSHI 6 6 500K
RBASSLO 6 9 500K

RVOLHI 7 3 1
RVOLLO 3 0 1MEG

RL 3 0 10MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END