* RC4558 OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* CREATED USING PARTS RELEASE 4.01 ON 09/08/89 AT 16:07
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | |
.SUBCKT RC4558   1 2 3 4 5
*
  C1   11 12 2.664E-12
  C2    6  7 20.00E-12
  DC    5 53 DX
  DE   54  5 DX
  DLP  90 91 DX
  DLN  92 90 DX
  DP    4  3 DX
  EGND 99  0 POLY(2) (3,0) (4,0) 0 .5 .5
  FB    7 99 POLY(5) VB VC VE VLP VLN 0 6.365E6 -6E6 6E6 6E6 -6E6
  GA 6  0 11 12 418.0E-6
  GCM   0  6 10 99 6.705E-9
  IEE   3 10 DC 34.28E-6
  HLIM 90  0 VLIM 1K
  Q1   11  2 13 QX
  Q2   12  1 14 QX
  R2    6  9 100.0E3
  RC1   4 11 2.652E3
  RC2   4 12 2.652E3
  RE1  13 10 1.122E3
  RE2  14 10 1.122E3
  REE  10 99 5.834E6
  RO1 8  5 125
  RO2 7 99 125
  RP    3  4 24.67E3
  VB    9  0 DC 0
  VC    3 53 DC 2.600
  VE   54  4 DC 2.600
  VLIM  7  8 DC 0
  VLP  91  0 DC 25
  VLN   0 92 DC 25
.MODEL DX D(IS=800.0E-18)
.MODEL QX PNP(IS=800.0E-18 BF=121.4)
.ENDS