Marshall classic three knob control

VIN 0 1 DC 0 AC 1
RS 1 2 1

C1 2 4 250P
R1 2 5 100K

RTREBLEHI 4 7 125K
RTREBLELO 7 6 125K

C2 5 6 100N
C3 5 9 47N

RMIDHI 9 9 5K
RMIDLO 9 0 5K

RBASSHI 6 6 125K
RBASSLO 6 9 125K

RVOLHI 7 3 1
RVOLLO 3 0 1MEG

RL 3 0 10MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END