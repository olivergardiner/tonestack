Marshall 18W single control

VIN 0 1 DC 0 AC 1
RS 1 2 47K

C1 2 4 10N

RTONELO 4 0 250K
RTONEHI 0 6 250K

R1 6 7 100K
C2 2 7 4.7N

RVOLHI 7 3 1
RVOLLO 3 0 1MEG

RL 3 0 1MEG

.OPTIONS NOACCT
.AC DEC 10 10 100K

.END